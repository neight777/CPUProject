library ieee;
use ieee.std_logic_1164.all;
entity SimpleCPU is
--Outputs you can display on fpga
port (
clk : in std_logic;
pcOut : out std_logic_vector(7 downto 0);
marOut : out std_logic_vector (7 downto 0);
irOutput : out std_logic_vector (7 downto 0);
mdriOutput : out std_logic_vector (7 downto 0);
mdroOutput : out std_logic_vector (7 downto 0);
aOut : out std_logic_vector (7 downto 0);
incrementOut : out std_logic
);
end;

architecture behavior of SimpleCPU is

signal pcRegOut  : std_logic_vector(7 downto 0);
signal marRegOut : std_logic_vector(7 downto 0);
signal mdroOut   : std_logic_vector(7 downto 0);
signal aRegOut   : std_logic_vector(7 downto 0);

--Initialize memory component
component memory_8_by_32
port( clk: in std_logic;
Write_Enable: in std_logic;
Read_Addr: in std_logic_vector (4 downto 0);
Data_in: in std_logic_vector (7 downto 0);
Data_out: out std_logic_vector(7 downto 0)
);
end component;

--initialize the alu
component ALU is
port(
  A     : in  std_logic_vector (7 downto 0);
  B     : in  std_logic_vector (7 downto 0);
  AluOp : in  std_logic_vector (2 downto 0);
  output: out std_logic_vector (7 downto 0)
);
end component;

--initialize the registers
component reg
port (
input : in std_logic_vector (7 downto 0);
output : out std_logic_vector (7 downto 0);
clk : in std_logic;
load : in std_logic
);
end component;

--initialize the program counter
component ProgramCounter
port (
increment : in std_logic;
clk : in std_logic;
output : out std_logic_vector (7 downto 0)
);
end component;

--initialize the mux
component TwoToOneMux
port (
A : in std_logic_vector (7 downto 0);
B : in std_logic_vector (7 downto 0);
address : in std_logic;
output : out std_logic_vector (7 downto 0)
);
end component;

--initialize the seven segment decoder
component sevenseg
port(
i : in std_logic_vector(3 downto 0);
o : out std_logic_vector(7 downto 0)
);
end component;

-- initialize control unit
component ControlUnit
port (
OpCode : in std_logic_vector(2 downto 0);
clk : in std_logic;
ToALoad : out std_logic;
ToMarLoad : out std_logic;
ToIrLoad : out std_logic;
ToMdriLoad : out std_logic;
ToMdroLoad : out std_logic;
ToPcIncrement : out std_logic;
ToMarMux : out std_logic;
ToRamWriteEnable : out std_logic;
ToAluOp : out std_logic_vector (2 downto 0)
);
end component;

-- Connections 
signal ramDataOutToMdri : std_logic_vector (7 downto 0);
-- MAR Multiplexer connections
signal pcToMarMux : std_logic_vector(7 downto 0);
signal muxToMar : std_logic_vector (7 downto 0);
-- RAM connections
signal marToRamReadAddr : std_logic_vector (4 downto 0);
signal mdroToRamDataIn : std_logic_vector (7 downto 0);
-- MDRI connections
signal mdriOut : std_logic_vector (7 downto 0);
-- IR connection
signal irOut : std_logic_vector (7 downto 0);
-- ALU / Accumulator connections
signal aluOut: std_logic_vector (7 downto 0);
signal aToAluB : std_logic_vector (7 downto 0);
-- Control Unit connections
signal cuToALoad : std_logic;
signal cuToMarLoad : std_logic;
signal cuToIrLoad : std_logic;
signal cuToMdriLoad : std_logic;
signal cuToMdroLoad : std_logic;
signal cuToPcIncrement : std_logic;
signal cuToMarMux : std_logic;
signal cuToRamWriteEnable : std_logic;
signal cuToAluOp : std_logic_vector (2 downto 0);
begin
--PORT MAP STATEMENTS
-- RAM
Map_Memory: memory_8_by_32 port map(clk=>clk,
Read_Addr=>marToRamReadAddr,
Data_in=>mdroToRamDataIn,
Data_Out=>ramDataOutToMdri,
Write_Enable=>cuToRamWriteEnable );

-- Accumulator
Map_A: reg port map(
  clk    => clk,
  load   => cuToALoad,
  input  => aluOut,
  output => aRegOut
);

-- ALU
MAP_ALU: ALU port map(
  A     => aToAluB,      
  B     => mdriOut,    
  AluOp => cuToAluOp,   
  output=> aluOut        
);


-- Program Counter
Map_PC: ProgramCounter port map(
  clk       => clk,
  increment => cuToPcIncrement,
  output    => pcRegOut
);


-- Instruction Register
Map_IR: reg port map(
  clk    => clk,
  load   => cuToIrLoad,
  input  => mdriOut,
  output => irOut
);


-- MAR mux
Map_MAR_Mux: TwoToOneMux port map(
  A       => pcRegOut,
  B       => irOut,
  address => cuToMarMux,
  output  => muxToMar
);

-- Memory Access Register
Map_MAR: reg port map(
  clk    => clk,
  load   => cuToMarLoad,
  input  => muxToMar,
  output => marRegOut
);


-- Memory Data Register Input
Map_MDRI: reg port map(clk=>clk,
input=>ramDataOutToMdri,
output=>mdriOut,
load=>cuToMdriLoad );


-- Memory Data Register Output
Map_MDRO: reg port map(
  clk    => clk,
  load   => cuToMdroLoad,
  input  => aRegOut,
  output => mdroOut
);




-- Control Unit
Map_CU: ControlUnit port map(
  OpCode          => irOut(7 downto 5),
  clk             => clk,
  ToALoad          => cuToALoad,
  ToMarLoad        => cuToMarLoad,
  ToIrLoad         => cuToIrLoad,
  ToMdriLoad       => cuToMdriLoad,
  ToMdroLoad       => cuToMdroLoad,
  ToPcIncrement    => cuToPcIncrement,
  ToMarMux         => cuToMarMux,
  ToRamWriteEnable => cuToRamWriteEnable,
  ToAluOp          => cuToAluOp
);

marToRamReadAddr <= marRegOut(4 downto 0);
mdroToRamDataIn  <= mdroOut;

pcOut        <= pcRegOut;
marOut       <= marRegOut;
irOutput     <= irOut;
mdriOutput   <= mdriOut;
mdroOutput   <= mdroOut;
aOut         <= aRegOut;
incrementOut <= cuToPcIncrement;


--would bind signals to fpga here but the cpu will be tested with the visual waveform tool
end behavior;